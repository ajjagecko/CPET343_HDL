-------------------------------------------------------------------------------
-- Andrew Akre
-- Structural Implementation of Single Bit Adder with Carry Over
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;     
use ieee.numeric_std.all; 

entity alu_and is
   port(
      a      :in std_logic;
      b      :in std_logic;
      x      :out std_logic;
   );
end alu_and;

architecture structural of alu_and is

begin

end